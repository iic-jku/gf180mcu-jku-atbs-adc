VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO gf180mcu_ws_ip__credits
  CLASS BLOCK ;
  FOREIGN gf180mcu_ws_ip__credits ;
  ORIGIN 0.000 0.000 ;
  SIZE 233.33 BY 100.0 ;
  OBS
      LAYER Metal5 ;
        RECT 0.0 0.0 233.33 100.0 ;
  END
END gf180mcu_ws_ip__credits
END LIBRARY