VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO gf180mcu_ws_ip__names
  CLASS BLOCK ;
  FOREIGN gf180mcu_ws_ip__names ;
  ORIGIN 0.000 0.000 ;
  SIZE 200.0 BY 200.0 ;
  OBS
      LAYER Metal5 ;
        RECT 0.0 0.0 200.0 200.0 ;
  END
END gf180mcu_ws_ip__names
END LIBRARY