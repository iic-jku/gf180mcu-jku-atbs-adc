library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.math_real.all;
package SpikesShiftRegSimVals is
--------------------------------------------------------
--SIMULATION CONSTANTS
--------------------------------------------------------
  constant CLK_FREQ: natural := 100000000;
  constant WIN_LENGTH: natural := 20;
  constant CNT_BITS : natural := 6;
  constant DATA_LENGTH : natural := 88;
  type T_SIM_SPIKES is array (0 to DATA_LENGTH - 1) of signed(CNT_BITS downto 0);
  constant SIM_SPIKES : T_SIM_SPIKES := (
"0011001", -- 25.000000 
"0100010", -- 34.000000 
"0101010", -- 42.000000 
"0110011", -- 51.000000 
"0111011", -- 59.000000 
"0000000", -- 0.000000 
"0000101", -- 5.000000 
"0001110", -- 14.000000 
"0011000", -- 24.000000 
"0100001", -- 33.000000 
"0101100", -- 44.000000 
"0110110", -- 54.000000 
"0000000", -- 0.000000 
"0000011", -- 3.000000 
"0001111", -- 15.000000 
"0011101", -- 29.000000 
"0101101", -- 45.000000 
"0000000", -- 0.000000 
"0000001", -- 1.000000 
"0011101", -- 29.000000 
"0000000", -- 0.000000 
"1000101", -- -59.000000 
"0000000", -- 0.000000 
"1110001", -- -15.000000 
"1100001", -- -31.000000 
"1010011", -- -45.000000 
"1000111", -- -57.000000 
"0000000", -- 0.000000 
"1111010", -- -6.000000 
"1110000", -- -16.000000 
"1100101", -- -27.000000 
"1011100", -- -36.000000 
"1010010", -- -46.000000 
"1001001", -- -55.000000 
"0000000", -- 0.000000 
"1111111", -- -1.000000 
"1110111", -- -9.000000 
"1101110", -- -18.000000 
"1100110", -- -26.000000 
"1011101", -- -35.000000 
"1010101", -- -43.000000 
"1001101", -- -51.000000 
"1000100", -- -60.000000 
"0000000", -- 0.000000 
"1111011", -- -5.000000 
"1110011", -- -13.000000 
"1101011", -- -21.000000 
"1100010", -- -30.000000 
"1011010", -- -38.000000 
"1010001", -- -47.000000 
"1001001", -- -55.000000 
"0000000", -- 0.000000 
"1111111", -- -1.000000 
"1110110", -- -10.000000 
"1101100", -- -20.000000 
"1100011", -- -29.000000 
"1011000", -- -40.000000 
"1001110", -- -50.000000 
"1000010", -- -62.000000 
"0000000", -- 0.000000 
"1110101", -- -11.000000 
"1100111", -- -25.000000 
"1010111", -- -41.000000 
"1000100", -- -60.000000 
"0000000", -- 0.000000 
"1100111", -- -25.000000 
"0000000", -- 0.000000 
"0110111", -- 55.000000 
"0000000", -- 0.000000 
"0001011", -- 11.000000 
"0011011", -- 27.000000 
"0101001", -- 41.000000 
"0110101", -- 53.000000 
"0000000", -- 0.000000 
"0000010", -- 2.000000 
"0001100", -- 12.000000 
"0010111", -- 23.000000 
"0100000", -- 32.000000 
"0101010", -- 42.000000 
"0110011", -- 51.000000 
"0111100", -- 60.000000 
"0000000", -- 0.000000 
"0000101", -- 5.000000 
"0001110", -- 14.000000 
"0010110", -- 22.000000 
"0011111", -- 31.000000 
"0100111", -- 39.000000 
"0101111");-- 47.000000 


end package SpikesShiftRegSimVals;
