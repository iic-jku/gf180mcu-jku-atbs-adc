library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package Spike2ThermoSimVals is

  constant THERMO_BITS: natural := 10;
  
end package Spike2ThermoSimVals;
