module gf180mcu_ws_ip__jku;
endmodule
