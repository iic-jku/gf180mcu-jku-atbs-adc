VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO gf180mcu_ws_ip__iicqc
  CLASS BLOCK ;
  FOREIGN gf180mcu_ws_ip__iicqc ;
  ORIGIN 0.000 0.000 ;
  SIZE 633.33 BY 100.0 ;
  OBS
      LAYER Metal5 ;
        RECT 0.0 0.0 633.33 100.0 ;
  END
END gf180mcu_ws_ip__iicqc
END LIBRARY